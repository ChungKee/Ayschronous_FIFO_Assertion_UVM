class AsynFIFO_sequence_item extends uvm_sequence_item;
    `uvm_object_utils(AsynFIFO_sequence_item)
    
    
  
    function new(string name = "AsynFIFO_sequence_item");
        super.new(name);
    endfunction
 
endclass : AsynFIFO_sequence_item